*
*
*
*                       LINUX           Fri Nov 14 00:11:38 2025
*
*
*
*  PROGRAM  advgen
*
*  Name           : advgen - Quantus QRC - (64-bit)
*  Version        : 15.2.7-s638
*  Build Date     : Wed Jan  4 18:11:53 PST 2017
*
*  HSPICE LIBRARY
*
*
*

*
.SUBCKT TSPCFF VDD! VSS! ck d q
*
*
*  caps2d version: 10
*
*
*       TRANSISTOR CARDS
*
*
MXinv_ck/Mmn0	ckb#11	ck#3	VSS!#14	VSS!#1	g45n1svt
+ L=4.5e-08	W=1.45e-07
+ AD=2.03e-14	AS=2.03e-14	PD=5.7e-07	PS=5.7e-07
+ NRD=3.388E-01	NRS=3.388E-01
+ scc=0.0026534 scb=0.0335332 sca=27.7828 sb=1.4e-07 sa=1.4e-07
Mmn1	a	d#3	VSS!#13	VSS!#1	g45n1svt	L=4.5e-08
+ W=1.45e-07
+ AD=8.7e-15	AS=8.7e-15	PD=4.9e-07	PS=4.9e-07
+ NRD=2.000E-01	NRS=3.388E-01
+ scc=0.000389368 scb=0.0118651 sca=11.7532 sb=2.45e-07 sa=1.4e-07
Mmn4	x#5	ckb#5	a	VSS!#1	g45n1svt	L=4.5e-08
+ W=1.45e-07
+ AD=2.03e-14	AS=2.03e-14	PD=4.9e-07	PS=4.9e-07
+ NRD=3.388E-01	NRS=2.000E-01
+ scc=0.000387736 scb=0.0112192 sca=11.1802 sb=1.4e-07 sa=2.45e-07
Mmn2	y#5	ckb	VSS!#12	VSS!#1	g45n1svt	L=4.5e-08
+ W=1.45e-07
+ AD=2.32e-14	AS=2.32e-14	PD=5.9e-07	PS=5.9e-07
+ NRD=3.388E-01	NRS=3.388E-01
+ scc=0.00038747 scb=0.0108541 sca=10.6844 sb=3.45e-07 sa=1.4e-07
Mmn3	qb#6	y#3	VSS!#12	VSS!#1	g45n1svt	L=4.5e-08
+ W=1.45e-07
+ AD=2.03e-14	AS=2.03e-14	PD=5.9e-07	PS=5.9e-07
+ NRD=3.388E-01	NRS=3.388E-01
+ scc=0.000387712 scb=0.0112005 sca=11.16 sb=1.4e-07 sa=3.45e-07
MXinv_q/Mmn0	q#1	qb#3	VSS!#11	VSS!#1	g45n1svt
+ L=4.5e-08	W=2.6e-07
+ AD=3.64e-14	AS=3.64e-14	PD=8e-07	PS=8e-07
+ NRD=2.046E-01	NRS=2.046E-01
+ scc=0.00232739 scb=0.0298965 sca=25.245 sb=1.4e-07 sa=1.4e-07
MXinv_ck/Mmp0	ckb#9	ck#1	VDD!#14	VDD!#1	g45p1svt
+ L=4.5e-08	W=2.15e-07
+ AD=3.01e-14	AS=3.01e-14	PD=7.1e-07	PS=7.1e-07
+ NRD=2.353E-01	NRS=2.353E-01
+ scc=0.00239434 scb=0.0309575 sca=27.6837 sb=1.4e-07 sa=1.4e-07
Mmp1	x#4	d#1	VDD!#10	VDD!#1	g45p1svt	L=4.5e-08
+ W=2.15e-07
+ AD=3.44e-14	AS=3.44e-14	PD=7.3e-07	PS=7.3e-07
+ NRD=2.353E-01	NRS=2.353E-01
+ scc=0.000130307 scb=0.00928939 sca=11.654 sb=4.5e-07 sa=1.4e-07
Mmp2	b	ckb#6	VDD!#10	VDD!#1	g45p1svt	L=4.5e-08
+ W=2.15e-07
+ AD=1.29e-14	AS=1.29e-14	PD=6.5e-07	PS=6.5e-07
+ NRD=1.349E-01	NRS=2.353E-01
+ scc=0.000128445 scb=0.00838672 sca=10.7652 sb=2.45e-07 sa=3.45e-07
Mmp4	y#6	x	b	VDD!#1	g45p1svt	L=4.5e-08
+ W=2.15e-07
+ AD=3.01e-14	AS=3.01e-14	PD=6.3e-07	PS=6.3e-07
+ NRD=2.353E-01	NRS=1.349E-01
+ scc=0.000128409 scb=0.00828104 sca=10.5904 sb=1.4e-07 sa=4.5e-07
Mmp3	c	y	VDD!#6	VDD!#1	g45p1svt	L=4.5e-08
+ W=2.15e-07
+ AD=1.29e-14	AS=1.29e-14	PD=6.3e-07	PS=6.3e-07
+ NRD=1.349E-01	NRS=2.353E-01
+ scc=0.000128651 scb=0.00862472 sca=11.0609 sb=2.45e-07 sa=1.4e-07
Mmp5	qb#4	ckb#7	c	VDD!#1	g45p1svt	L=4.5e-08
+ W=2.15e-07
+ AD=3.01e-14	AS=3.01e-14	PD=6.3e-07	PS=6.3e-07
+ NRD=2.353E-01	NRS=1.349E-01
+ scc=0.000130139 scb=0.00924431 sca=11.619 sb=1.4e-07 sa=2.45e-07
MXinv_q/Mmp0	q#2	qb	VDD!#3	VDD!#1	g45p1svt	L=4.5e-08
+ W=3.9e-07
+ AD=5.46e-14	AS=5.46e-14	PD=1.06e-06	PS=1.06e-06
+ NRD=1.364E-01	NRS=1.364E-01
+ scc=0.00229311 scb=0.0313093 sca=27.4572 sb=1.4e-07 sa=1.4e-07
*
*
*       RESISTOR AND CAP/DIODE CARDS
*
Rl1	ck#1	ck#2	  173.7687
Rl2	ck#2	ck#3	  158.3841
Rl3	d#1	d#2	  129.5379
Rl4	d#2	d#3	  202.6149
Rl5	x	x#2	  115.3867
Rl6	ckb	ckb#2	  138.2566
Rl7	ckb#2	ckb#3	  111.9279
Rl8	ckb#3	ckb#4	   11.9279
Rl9	ckb#4	ckb#5	  138.2566
Rl10	ckb#3	ckb#6	  180.4507
Rl11	y	y#2	  116.5405
Rl12	y#2	y#3	  212.6944
Rl13	ckb#7	ckb#8	  211.0764
Rl14	qb	qb#2	  106.4610
Rl15	qb#2	qb#3	  114.1533
Rk1	ck#2	ck	   45.0552
Rk2	d#2	d	   45.0572
Rk3	ckb#9	ckb#10	   62.4819
Rk4	ckb#10	ckb#11	   75.3353
Rk5	ckb#10	ckb#4	   45.2960
Rk6	x#2	x#3	5.119E-02
Rk7	x#3	x#4	   62.5383
Rk8	x#3	x#5	   75.6540
Rk9	y#2	y#4	   45.1281
Rk10	y#4	y#5	   75.6160
Rk11	y#4	y#6	   62.3725
Rk12	ckb#2	ckb#8	   45.2162
Rk13	qb#4	qb#5	   62.4807
Rk14	qb#5	qb#6	   75.4759
Rk15	qb#5	qb#2	   45.1205
Rk16	q	q#1	   37.8260
Rk17	q	q#2	   21.0277
Rk18	VDD!#1	VDD!#2	   75.1110
Rk19	VDD!#2	VDD!#3	   20.9649
Rk20	VDD!#2	VDD!#4	    0.1104
Rk21	VDD!#4	VDD!#5	    0.1104
Rk22	VDD!#5	VDD!#6	   62.2128
Rk23	VDD!#5	VDD!#7	    0.1110
Rk24	VDD!#7	VDD!#8	    0.1129
Rk25	VDD!#8	VDD!#9	4.748E-02
Rk26	VDD!#9	VDD!#10	   62.1999
Rk27	VDD!#9	VDD!#11	6.505E-02
Rk28	VDD!#11	VDD!#12	    0.1129
Rk29	VDD!#12	VDD!	    0.1129
Rk31	VDD!	VDD!#14	   62.2240
Rk32	VDD!#1	VDD!#2	   75.0000
Rk33	VDD!#1	VDD!#4	   75.0000
Rk34	VDD!#1	VDD!#5	   75.0000
Rk35	VDD!#1	VDD!#7	   75.0000
Rk36	VDD!#1	VDD!#8	   75.0000
Rk37	VDD!#1	VDD!#11	   75.0000
Rk38	VDD!#1	VDD!#12	   75.0000
Rk39	VDD!#1	VDD!	   75.0000
Rk40	VSS!#1	VSS!#2	   62.1110
Rk41	VSS!#2	VSS!#3	    0.1104
Rk42	VSS!#3	VSS!#4	    0.1104
Rk43	VSS!#4	VSS!#5	    0.1110
Rk44	VSS!#5	VSS!#6	    0.1129
Rk45	VSS!#6	VSS!#7	    0.1129
Rk46	VSS!#7	VSS!#8	3.745E-02
Rk47	VSS!#8	VSS!#9	7.509E-02
Rk48	VSS!#9	VSS!	    0.1129
Rk50	VSS!#2	VSS!#11	   37.7315
Rk51	VSS!#4	VSS!#12	   75.1974
Rk52	VSS!#8	VSS!#13	   75.1775
Rk53	VSS!	VSS!#14	   75.2016
Rk54	VSS!#1	VSS!#2	   62.0000
Rk55	VSS!#1	VSS!#3	   62.0000
Rk56	VSS!#1	VSS!#4	   62.0000
Rk57	VSS!#1	VSS!#5	   62.0000
Rk58	VSS!#1	VSS!#6	   62.0000
Rk59	VSS!#1	VSS!#7	   62.0000
Rk60	VSS!#1	VSS!#9	   62.0000
Rk61	VSS!#1	VSS!	   62.0000
*
*       CAPACITOR CARDS
*
*
C1	ckb#3	y#2	3.09493E-18
C2	ck	VDD!	2.01491E-19
C3	VSS!#1	q#1	7.97298E-18
C4	ckb#5	VDD!#1	6.98069E-18
C5	y#4	VDD!#6	2.22051E-18
C6	ckb#9	d#1	1.22472E-18
C7	ckb#2	y#2	2.48786E-17
C8	x#5	ckb#4	2.9573E-18
C9	VDD!	d#1	3.49167E-19
C10	VDD!	ck#1	5.40627E-18
C11	VDD!#10	ck#1	2.02294E-19
C12	y#4	ckb#8	2.54129E-18
C13	x#3	y#6	9.31046E-18
C14	ck#2	VDD!	7.41989E-19
C15	x#2	y#2	3.94958E-18
C16	d#3	VDD!#1	9.72236E-18
C17	y#6	VDD!#6	1.90509E-17
C18	q#1	VDD!#1	6.62528E-18
C19	VSS!#1	ck#3	1.7878E-19
C20	qb#5	ckb#8	4.78201E-17
C21	qb#5	ckb#7	5.37569E-19
C22	x#3	y#2	4.90883E-19
C23	ckb#9	ck#1	5.83862E-18
C24	VSS!#12	qb#6	1.35282E-17
C25	x#5	d#2	3.24791E-19
C26	VSS!#1	qb#6	7.30903E-18
C27	ckb#2	x#2	3.00082E-18
C28	VDD!#14	ck#1	2.99015E-18
C29	ck#3	VDD!#1	1.58537E-17
C30	VSS!#13	ckb#4	1.61419E-18
C31	VSS!#11	VDD!#1	1.58585E-18
C32	VSS!#1	qb#2	2.36564E-18
C33	ck	VDD!#1	8.52365E-18
C34	y#5	qb#6	6.7325E-18
C35	qb#2	VDD!#1	1.59052E-17
C36	y#2	qb#5	1.04442E-17
C37	ckb#3	x#2	1.0762E-17
C38	VSS!#1	ckb#8	2.46549E-18
C39	qb#6	VDD!#1	3.18045E-18
C40	qb#2	q	3.12627E-17
C41	d	ck#2	6.53112E-19
C42	ck	VDD!#14	1.95394E-18
C43	VSS!#1	y#5	7.42275E-18
C44	d	VDD!#1	4.08976E-18
C45	q#1	qb#3	5.57259E-18
C46	x#3	VDD!#10	6.50798E-18
C47	y#4	ckb#2	3.75278E-17
C48	ckb#8	VDD!#1	1.5011E-17
C49	VSS!#12	VDD!#1	4.97306E-19
C50	y#5	VSS!#12	1.35282E-17
C51	ckb#10	x#4	3.39721E-18
C52	VSS!#11	qb#3	3.99549E-18
C53	qb#2	VDD!#3	5.3766E-18
C54	VSS!#14	ck	2.07872E-18
C55	VDD!#10	y#6	1.28606E-17
C56	VSS!#1	x#5	1.25233E-17
C57	ckb#2	qb#5	1.97063E-18
C58	q	VDD!#1	1.46421E-17
C59	x#3	ckb#3	4.98705E-18
C60	d	x#4	3.1649E-18
C61	ckb#7	qb	6.32643E-18
C62	y#2	VDD!#1	1.26074E-17
C63	VSS!#1	ckb#2	3.43704E-18
C64	y#5	VDD!#1	3.32323E-18
C65	ckb#4	d#2	3.75805E-17
C66	VSS!#12	qb#3	2.5179E-19
C67	y#4	x#2	1.70077E-18
C68	x#3	ckb#6	1.83546E-18
C69	x#4	y#6	4.10208E-18
C70	y	ckb#7	4.13894E-17
C71	VSS!#11	y#3	1.40061E-18
C72	ckb#2	VDD!#1	1.15706E-17
C73	ckb#4	ck#2	2.07562E-19
C74	x#5	VDD!#1	5.27269E-18
C75	d#2	ckb#3	1.32656E-17
C76	qb#6	y#3	3.77638E-18
C77	ckb#10	d	2.51035E-17
C78	ckb#10	x#3	1.55051E-18
C79	ckb#4	x#3	2.40661E-17
C80	x	y	4.1989E-18
C81	VSS!#12	y#3	1.84043E-18
C82	x#2	VDD!#1	6.4307E-18
C83	VSS!#14	ck#2	3.3987E-18
C84	VSS!#1	ckb#4	5.17578E-18
C85	ck#2	d#2	9.65041E-18
C86	x#5	y#5	4.14478E-17
C87	ckb#10	d#2	6.14969E-18
C88	ckb#6	x	3.55652E-17
C89	VSS!#1	ckb#11	4.83211E-18
C90	qb#6	ckb	1.04389E-18
C91	ckb#4	VDD!#1	8.68397E-18
C92	x#3	d#2	1.51848E-17
C93	VSS!#13	VDD!#1	8.66372E-19
C94	x#4	VDD!#10	1.58073E-17
C95	VSS!#12	ckb	1.53267E-18
C96	VSS!#8	VDD!#1	2.31692E-18
C97	qb#5	q	1.01543E-17
C98	d#1	ckb#6	1.69542E-17
C99	ck#2	ckb#10	3.5609E-17
C100	y#2	VDD!#6	4.09409E-18
C101	d#2	VDD!#1	1.73491E-17
C102	y#5	ckb	3.05593E-18
C103	VSS!#8	ck#3	1.17207E-18
C104	ckb#11	VDD!#1	4.21749E-18
C105	VDD!#9	ckb#6	9.23033E-19
C106	ck#1	d#1	6.22494E-18
C107	VSS!#1	ckb#3	6.55623E-19
C108	x#5	ckb	1.09652E-18
C109	ckb#8	qb	1.73241E-18
C110	x#3	y#4	5.26857E-17
C111	ck#2	VDD!#1	2.61402E-17
C112	VDD!#6	ckb#2	7.17698E-19
C113	VSS!#14	VDD!#1	2.31691E-18
C114	y#5	ckb#5	1.09652E-18
C115	VSS!#1	ckb#10	1.46543E-18
C116	ckb#9	x#4	3.22334E-17
C117	VSS!#13	ckb	2.82157E-19
C118	y#6	ckb#2	5.84432E-19
C119	y#2	ckb#7	6.43305E-18
C120	VSS!#1	VDD!#1	3.93865E-18
C121	x#5	ckb#5	3.30939E-18
C122	ckb#3	VDD!#1	9.56142E-18
C123	VDD!#9	d#1	8.88403E-19
C124	VSS!#13	x#5	9.78812E-18
C125	y#3	qb#3	4.58839E-18
C126	y#6	x#2	2.23963E-18
C127	ckb#10	VDD!#1	1.39477E-17
C128	VSS!#13	ckb#5	5.81189E-19
C129	VSS!#1	y#4	5.70133E-19
C130	x#2	y	1.057E-18
C131	x#5	d#3	1.2238E-18
C132	VSS!#11	qb#2	5.02731E-18
C133	qb	VDD!#1	1.73397E-17
C134	ckb	y#3	1.61953E-17
C135	q#2	VDD!#1	1.38962E-17
C136	q#2	qb	5.60806E-18
C137	ckb#11	x#5	4.17362E-18
C138	x#3	VDD!#1	1.26284E-17
C139	y#4	qb#5	7.5119E-18
C140	VDD!#9	ck#1	4.72019E-19
C141	qb#5	q#1	1.30039E-18
C142	VDD!#14	ckb#9	1.86747E-17
C143	VSS!#1	qb#5	5.17723E-18
C144	VDD!#3	qb	5.27041E-18
C145	qb#5	y#3	7.43245E-19
C146	ckb#7	VDD!#1	1.01835E-17
C147	y#4	VDD!#1	9.52291E-18
C148	ckb#6	x#2	1.55194E-17
C149	VDD!#3	ckb#7	1.80961E-18
C150	VDD!#6	qb	4.05939E-19
C151	ckb#11	d#3	2.51624E-18
C152	y	VDD!#1	1.12001E-17
C153	qb#4	ckb#7	3.38257E-18
C154	qb#4	VDD!#1	9.56433E-18
C155	VDD!#3	q#2	3.15412E-17
C156	qb#5	VDD!#1	1.39544E-17
C157	d#2	ckb#6	3.43044E-18
C158	d#3	ckb#5	3.93734E-17
C159	VSS!#13	ck#3	1.52634E-18
C160	VDD!#6	ckb#7	6.95521E-19
C161	x	VDD!#1	8.85655E-18
C162	qb#4	y	9.3364E-19
C163	x#5	ckb#3	8.93514E-19
C164	ckb#11	ck#3	4.93764E-18
C165	ckb#11	VSS!#13	1.38007E-17
C166	ckb#10	d#3	1.04564E-18
C167	ckb#6	VDD!#1	9.99289E-18
C168	VDD!#6	y	2.47792E-18
C169	ck#3	d#3	5.88809E-18
C170	qb#5	q#2	5.67363E-18
C171	VSS!#12	y#2	8.195E-19
C172	VSS!#14	ck#3	2.51202E-18
C173	ck#1	d#2	1.02164E-18
C174	qb#4	VDD!#3	2.84868E-17
C175	ckb#2	y#3	4.49031E-18
C176	d#2	x#4	1.07855E-17
C177	ckb#10	x#5	4.52337E-18
C178	d#1	VDD!#1	1.07169E-17
C179	y#6	VDD!#1	9.58053E-18
C180	VDD!#6	x	1.06573E-18
C181	ckb#10	ck#3	5.47642E-19
C182	VSS!#12	ckb#2	4.76175E-18
C183	y#6	x	3.08452E-18
C184	VSS!#11	q#1	2.19832E-17
C185	qb#5	VDD!#3	4.32791E-18
C186	ck#1	VDD!#1	1.57629E-17
C187	VSS!#1	qb#3	5.68931E-18
C188	y#5	ckb#2	1.08708E-18
C189	y#4	qb#4	4.27213E-18
C190	VDD!#10	x	6.95521E-19
C191	VSS!#14	ckb#11	1.35282E-17
C192	y#6	ckb#6	1.13696E-18
C193	qb#3	VDD!#1	1.34761E-17
C194	ckb#8	qb#2	6.83785E-18
C195	qb#6	q#1	2.4756E-18
C196	VSS!#1	y#3	5.29024E-18
C197	y#5	qb#5	2.26489E-18
C198	ck#2	VDD!#14	3.20555E-18
C199	VDD!#6	qb#4	1.28606E-17
C200	y#2	qb#2	2.18628E-18
C201	x#5	y#4	7.57631E-18
C202	VDD!#10	ckb#6	2.02918E-18
C203	y#3	VDD!#1	1.0484E-17
C204	VSS!#13	ckb#10	2.73768E-18
C205	x#4	VDD!#1	7.74152E-18
C206	d#3	ckb#4	8.00209E-18
C207	VSS!#1	ckb	3.67207E-18
C208	x#4	ckb#6	1.07095E-18
C209	ckb#8	y#2	4.43115E-17
C210	qb#6	VSS!#11	1.61157E-17
C211	y#6	qb#4	1.14619E-18
C212	ckb	VDD!#1	7.69041E-18
C213	VDD!#10	d#1	1.7468E-18
C214	ckb#9	VDD!#1	1.24796E-17
C215	y#4	qb	7.75514E-19
C216	VSS!#1	ckb#5	2.4886E-18
C217	x#4	d#1	3.15618E-18
C218	ck#2	d#3	1.02339E-18
C219	y#3	qb#2	1.74487E-19
C220	y#5	qb#3	2.821E-19
C221	VDD!#10	y	2.95047E-19
C222	VDD!#10	ckb#4	6.34144E-19
C223	VSS!#12	ckb#5	1.73807E-19
C224	VSS!#8	ckb	1.86344E-19
C225	VSS!#8	ckb#5	2.21461E-19
C226	qb#5	ckb#4	2.45418E-19
C227	qb#6	ckb#5	3.14064E-19
C228	x#4	y#4	2.31066E-19
C229	y#4	ckb#4	2.71358E-19
C230	y#4	ckb#3	3.32741E-19
C231	y#4	ckb#7	4.75371E-19
C232	q#1	qb#2	1.43615E-19
C233	x#3	ckb#2	3.35849E-19
C234	VDD!	VSS!	1.379E-19
C235	ck	VSS!	2.33329E-19
C236	q	VSS!	4.94013E-19
C237	a	VSS!	2.73015E-19
C238	c	VSS!	4.47876E-19
C239	b	VSS!	4.47876E-19
C240	qb	VSS!	1.20852E-19
C241	ckb#7	VSS!	4.23428E-19
C242	y	VSS!	7.57858E-19
C243	x	VSS!	9.10916E-19
C244	ckb#6	VSS!	5.25346E-19
C245	d#1	VSS!	1.10841E-18
C246	ck#1	VSS!	2.75051E-18
C247	y#3	VSS!	6.51725E-19
C248	ckb	VSS!	1.1892E-19
C249	ckb#5	VSS!	1.36508E-19
C250	d#3	VSS!	7.25793E-18
C251	ck#3	VSS!	6.15777E-18
C252	qb#2	VSS!	2.32862E-19
C253	ckb#8	VSS!	6.553E-19
C254	y#2	VSS!	5.9501E-19
C255	ckb#2	VSS!	4.3617E-19
C256	x#2	VSS!	6.92496E-19
C257	ckb#4	VSS!	2.00375E-19
C258	d#2	VSS!	1.15113E-18
C259	ck#2	VSS!	2.71658E-18
C260	VDD!#1	VSS!	3.40184E-18
C261	q#2	VSS!	5.27315E-19
C262	VDD!#3	VSS!	2.26745E-19
C263	qb#4	VSS!	4.86235E-19
C264	VDD!#6	VSS!	1.33079E-19
C265	y#6	VSS!	1.47479E-18
C266	x#4	VSS!	2.86223E-18
C267	ckb#9	VSS!	1.73427E-19
C268	VDD!#14	VSS!	2.08743E-19
C269	q#1	VSS!	4.90969E-19
C270	qb#6	VSS!	1.8348E-19
C271	y#5	VSS!	1.7657E-19
C272	x#5	VSS!	1.82541E-18
C273	ckb#3	VSS!	7.69356E-21
C274	ckb#10	VSS!	3.74053E-19
C275	x#3	VSS!	1.47373E-19
C276	y#4	VSS!	1.40081E-19
C277	qb#5	VSS!	4.32259E-19
C278	VDD!#9	VSS!	4.81665E-19
*
*
.ENDS TSPCFF
*
